`ifndef PROGRAM_VH
`define PROGRAM_VH

DATA_MEMORY(0,  LDI, -11'd4};
DATA_MEMORY(1,  STO,  11'd1};
DATA_MEMORY(2,  LDI,  11'd2};
DATA_MEMORY(3,  ADD,  11'd1};
DATA_MEMORY(4,  STO,  11'd2};
DATA_MEMORY(5,  LDI,  11'd123};
DATA_MEMORY(6,  ADDI, 11'd7 };
DATA_MEMORY(7,  LD,   11'd2};
DATA_MEMORY(8,  ADDI  11'd4};
DATA_MEMORY(9,  SUBI  11'd50};
DATA_MEMORY(10, SUB,  11'd1};
DATA_MEMORY(11, HLT,  11'd0};

`undef DATA_MEMORY

`endif



