`ifndef CONSTANTS_VH
`define CONSTANTS_VH

`define PROC_BITS 32        // General processor bit size
`define REG_ADDRS_BITS 5    // Registers addresses bit size
`define PC_BITS 8
`define OPCODE_BITS 6
`define INSTRUCTION_BITS 32

`endif
