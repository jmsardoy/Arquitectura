`ifndef INSTRUCTIONS_VH
`define INSTRUCTIONS_VH

INSTRUCTION(HLT, 'b00000)
INSTRUCTION(STO, 'b00001)
INSTRUCTION(LD,  'b00010)
INSTRUCTION(LDI, 'b00011)
INSTRUCTION(ADD, 'b00100)
INSTRUCTION(ADDI,'b00101)
INSTRUCTION(SUB, 'b00110)
INSTRUCTION(SUBI,'b00111)

`undef `INSTRUCTION

`endif
