`ifndef MEMORY_DEFS_VH
`define MEMORY_DEFS_VH

`define ADDRESS_BITS 11
`define DATA_BITS 16

`endif
